-- fadfaf